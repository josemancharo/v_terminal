module commands
import app_state {Command, AppState}
import types { Primitive }

pub fn define_function(mut state &AppState, params []string) Primitive {
	return 0
}