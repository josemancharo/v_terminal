module types

pub union Primitive {
	int
	string
	bool
	f32
}