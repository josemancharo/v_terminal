module types

pub struct Function {
	pub:
		params []string
		definition string
}