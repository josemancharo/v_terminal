module util

pub fn parse_parameters(params []string){

}